module pipelined_computer (clock,btn,sw,seven,vga_r,vga_g,vga_b,clk_vga,hsync,vsync,VGA_BLANK_N,VGA_SYNC_N);
	input clock,btn;
   input [17:0] sw;
   
   output [55:0] seven;
   output [9:0] vga_r,vga_g,vga_b;
   output clk_vga,hsync,vsync,VGA_BLANK_N,VGA_SYNC_N;

	wire resetn;
	wire [31:0] in_port0,in_port1,in_port2;
	wire [31:0] out_port0,out_port1,out_port2;
	wire [31:0] pc,ealu,malu,walu;
	
	wire [31:0] bpc,jpc,npc,pc4,ins, inst;
	wire [31:0] dpc4,da,db,dimm;
	wire [31:0] epc4,ea,eb,eimm;
	wire [31:0] mb,mmo;
	wire [31:0] wmo,wdi;
	wire [4:0] drn,ern0,ern,mrn,wrn;
	wire [3:0] daluc,ealuc;
	wire [1:0] pcsource;
	wire wpcir;
	wire dwreg,dm2reg,dwmem,daluimm,dshift,djal;
	wire ewreg,em2reg,ewmem,ealuimm,eshift,ejal;
	wire mwreg,mm2reg,mwmem;
	wire wwreg,wm2reg;
	wire mem_clock = ~clock;
	
	assign in_port0[7:0] = sw[7:0];
	assign in_port0[31:8] = 24'b0;
	assign in_port1[7:0] = sw[15:8];
	assign in_port1[31:8] = 24'b0;
	assign in_port2[1:0] = sw[17:16];
	assign in_port2[31:2] = 24'b0;
	assign resetn = btn;
	
	digit seven_dig(out_port1[7:0], out_port0[7:0], out_port2[7:0], seven[55:0]);
	vga_display vga_d(clock,resetn,in_port2[1:0],out_port1[7:0],out_port0[7:0],out_port2[7:0],vga_r,vga_g,vga_b,clk_vga,hsync,vsync,VGA_BLANK_N,VGA_SYNC_N);
	
	pipepc prog_cnt (npc,wpcir,clock,resetn,pc);
	pipeif if_stage (pcsource,pc,bpc,da,jpc,npc,pc4,ins,mem_clock);
	pipeir inst_reg (pc4,ins,wpcir,clock,resetn,dpc4,inst);
	pipeid id_stage (mwreg,mrn,ern,ewreg,em2reg,mm2reg,dpc4,inst,
	wrn,wdi,ealu,malu,mmo,wwreg,clock,resetn,
	bpc,jpc,pcsource,wpcir,dwreg,dm2reg,dwmem,daluc,
	daluimm,da,db,dimm,drn,dshift,djal);
	pipedereg de_reg (dwreg,dm2reg,dwmem,daluc,daluimm,da,db,dimm,drn,dshift,
	djal,dpc4,clock,resetn,ewreg,em2reg,ewmem,ealuc,ealuimm,
	ea,eb,eimm,ern0,eshift,ejal,epc4);
	pipeexe exe_stage (ealuc,ealuimm,ea,eb,eimm,eshift,ern0,epc4,ejal,ern,ealu);
	pipeemreg em_reg (ewreg,em2reg,ewmem,ealu,eb,ern,clock,resetn,
	mwreg,mm2reg,mwmem,malu,mb,mrn);
	pipemem mem_stage (mwmem,malu,mb,clock,mem_clock,mmo,resetn,in_port0,in_port1,in_port2,out_port0,out_port1,out_port2);
	pipemwreg mw_reg (mwreg,mm2reg,mmo,malu,mrn,clock,resetn,
	wwreg,wm2reg,wmo,walu,wrn);
	mux2x32 wb_stage (walu,wmo,wm2reg,wdi);
endmodule
